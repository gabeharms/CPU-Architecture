`timescale 1ns / 1ps
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//
// Author      : Gabe Harms
// Create Date : 03/20/12	
// Module Name : Sign Extention    
// Project Name: CPU_Datapath
//
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

module instruction_memory

(
	address,
	instruction
);

    //--------------------------
	// Parameters
	//--------------------------	
	
    //--------------------------
	// Input Ports
	//--------------------------
	// < Enter Input Ports  >
	input		[31:0]	address;
	
    //--------------------------
    // Output Ports
    //--------------------------
    // < Enter Output Ports  >	
    output 	reg [31:0] 	instruction;
		
    //--------------------------
    // Bidirectional Ports
    //--------------------------
    // < Enter Bidirectional Ports in Alphabetical Order >
    // None
      
    ///////////////////////////////////////////////////////////////////
    // Begin Design
    ///////////////////////////////////////////////////////////////////
    //-------------------------------------------------
    // Signal Declarations: local params
    //-------------------------------------------------
   
    //-------------------------------------------------
    // Signal Declarations: reg
    //-------------------------------------------------    
    reg	[31:0] instruction_memory	[255:0];
	
    //-------------------------------------------------
    // Signal Declarations: wire
    //-------------------------------------------------
		
	//---------------------------------------------------------------
	// Instantiations
	//---------------------------------------------------------------
	// None

	//---------------------------------------------------------------
	// Combinatorial Logic
	//---------------------------------------------------------------
	initial
	begin
		$readmemh("program.mips",instruction_memory);
	end
	
	always @ ( * )
	begin
	instruction = instruction_memory[address[9:2]];
	end
	
 endmodule  



